`define sil   32'd50000000 // slience

module music_L_ch (
	input [9:0] ibeatNum,
	input state_for_L_ch,
	output reg [31:0] toneL,
    output reg [31:0] toneR
);
/*--------------------------------*/
//↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓↓
//For state_for_L_ch
//parameter 
//  waiting_deposit = 1'b0,
//  waiting_playing = 1'b1;
//For state_for_L_ch
//↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑↑
/*--------------------------------*/

    always @* begin
        toneR = `sil;
    end

    always @(*) begin
        if (state_for_L_ch == 1'b0/*waiting_deposit*/) begin
            case(ibeatNum)
                12'd0: toneL = 32'd524; 12'd1: toneL = 32'd524; 
                12'd2: toneL = 32'd524; 12'd3: toneL = `sil; 
                12'd4: toneL = 32'd698; 12'd5: toneL = 32'd698; 
                12'd6: toneL = 32'd698; 12'd7: toneL = `sil; 
                12'd8: toneL = 32'd880; 12'd9: toneL = 32'd880; 
                12'd10: toneL = 32'd880; 12'd11: toneL = `sil; 
                12'd12: toneL = 32'd1048; 12'd13: toneL = 32'd1048; 
                12'd14: toneL = 32'd1048; 12'd15: toneL = `sil; 
                12'd16: toneL = 32'd1048; 12'd17: toneL = 32'd1048; 
                12'd18: toneL = 32'd1048; 12'd19: toneL = `sil; 
                12'd20: toneL = 32'd1396; 12'd21: toneL = 32'd1396; 
                12'd22: toneL = 32'd1396; 12'd23: toneL = `sil; 
                12'd24: toneL = 32'd1760; 12'd25: toneL = 32'd1760; 
                12'd26: toneL = 32'd1760; 12'd27: toneL = `sil; 
                12'd28: toneL = 32'd2096; 12'd29: toneL = 32'd2096; 
                12'd30: toneL = 32'd2096; 12'd31: toneL = `sil; 
                12'd32: toneL = 32'd2096; 12'd33: toneL = 32'd2096; 
                12'd34: toneL = 32'd2096; 12'd35: toneL = `sil; 
                12'd36: toneL = 32'd1760; 12'd37: toneL = 32'd1760; 
                12'd38: toneL = 32'd1760; 12'd39: toneL = `sil; 
                12'd40: toneL = 32'd1396; 12'd41: toneL = 32'd1396; 
                12'd42: toneL = 32'd1396; 12'd43: toneL = `sil; 
                12'd44: toneL = 32'd1048; 12'd45: toneL = 32'd1048; 
                12'd46: toneL = 32'd1048; 12'd47: toneL = `sil; 
                12'd48: toneL = 32'd1048; 12'd49: toneL = 32'd1048; 
                12'd50: toneL = 32'd1048; 12'd51: toneL = `sil; 
                12'd52: toneL = 32'd880; 12'd53: toneL = 32'd880; 
                12'd54: toneL = 32'd880; 12'd55: toneL = `sil; 
                12'd56: toneL = 32'd698; 12'd57: toneL = 32'd698; 
                12'd58: toneL = 32'd698; 12'd59: toneL = `sil; 
                12'd60: toneL = 32'd524; 12'd61: toneL = 32'd524; 
                12'd62: toneL = 32'd524; 12'd63: toneL = `sil; 
                12'd64: toneL = 32'd524; 12'd65: toneL = 32'd524; 
                12'd66: toneL = 32'd524; 12'd67: toneL = `sil; 
                12'd68: toneL = 32'd660; 12'd69: toneL = 32'd660; 
                12'd70: toneL = 32'd660; 12'd71: toneL = `sil; 
                12'd72: toneL = 32'd784; 12'd73: toneL = 32'd784; 
                12'd74: toneL = 32'd784; 12'd75: toneL = `sil; 
                12'd76: toneL = 32'd1048; 12'd77: toneL = 32'd1048; 
                12'd78: toneL = 32'd1048; 12'd79: toneL = `sil; 
                12'd80: toneL = 32'd1048; 12'd81: toneL = 32'd1048; 
                12'd82: toneL = 32'd1048; 12'd83: toneL = `sil; 
                12'd84: toneL = 32'd1320; 12'd85: toneL = 32'd1320; 
                12'd86: toneL = 32'd1320; 12'd87: toneL = `sil; 
                12'd88: toneL = 32'd1568; 12'd89: toneL = 32'd1568; 
                12'd90: toneL = 32'd1568; 12'd91: toneL = `sil; 
                12'd92: toneL = 32'd2096; 12'd93: toneL = 32'd2096; 
                12'd94: toneL = 32'd2096; 12'd95: toneL = `sil; 
                12'd96: toneL = 32'd2096; 12'd97: toneL = 32'd2096; 
                12'd98: toneL = 32'd2096; 12'd99: toneL = `sil; 
                12'd100: toneL = 32'd1568; 12'd101: toneL = 32'd1568; 
                12'd102: toneL = 32'd1568; 12'd103: toneL = `sil; 
                12'd104: toneL = 32'd1320; 12'd105: toneL = 32'd1320; 
                12'd106: toneL = 32'd1320; 12'd107: toneL = `sil; 
                12'd108: toneL = 32'd1048; 12'd109: toneL = 32'd1048; 
                12'd110: toneL = 32'd1048; 12'd111: toneL = `sil; 
                12'd112: toneL = 32'd1048; 12'd113: toneL = 32'd1048; 
                12'd114: toneL = 32'd1048; 12'd115: toneL = `sil; 
                12'd116: toneL = 32'd784; 12'd117: toneL = 32'd784; 
                12'd118: toneL = 32'd784; 12'd119: toneL = `sil; 
                12'd120: toneL = 32'd660; 12'd121: toneL = 32'd660; 
                12'd122: toneL = 32'd660; 12'd123: toneL = `sil; 
                12'd124: toneL = 32'd524; 12'd125: toneL = 32'd524; 
                12'd126: toneL = 32'd524; 12'd127: toneL = `sil; 
                12'd128: toneL = 32'd588; 12'd129: toneL = 32'd588; 
                12'd130: toneL = 32'd588; 12'd131: toneL = `sil; 
                12'd132: toneL = 32'd698; 12'd133: toneL = 32'd698; 
                12'd134: toneL = 32'd698; 12'd135: toneL = `sil; 
                12'd136: toneL = 32'd880; 12'd137: toneL = 32'd880; 
                12'd138: toneL = 32'd880; 12'd139: toneL = `sil; 
                12'd140: toneL = 32'd1048; 12'd141: toneL = 32'd1048; 
                12'd142: toneL = 32'd1048; 12'd143: toneL = `sil; 
                12'd144: toneL = 32'd1176; 12'd145: toneL = 32'd1176; 
                12'd146: toneL = 32'd1176; 12'd147: toneL = `sil; 
                12'd148: toneL = 32'd1396; 12'd149: toneL = 32'd1396; 
                12'd150: toneL = 32'd1396; 12'd151: toneL = `sil; 
                12'd152: toneL = 32'd1760; 12'd153: toneL = 32'd1760; 
                12'd154: toneL = 32'd1760; 12'd155: toneL = `sil; 
                12'd156: toneL = 32'd2096; 12'd157: toneL = 32'd2096; 
                12'd158: toneL = 32'd2096; 12'd159: toneL = `sil; 
                12'd160: toneL = 32'd2096; 12'd161: toneL = 32'd2096; 
                12'd162: toneL = 32'd2096; 12'd163: toneL = `sil; 
                12'd164: toneL = 32'd1760; 12'd165: toneL = 32'd1760; 
                12'd166: toneL = 32'd1760; 12'd167: toneL = `sil; 
                12'd168: toneL = 32'd1396; 12'd169: toneL = 32'd1396; 
                12'd170: toneL = 32'd1396; 12'd171: toneL = `sil; 
                12'd172: toneL = 32'd1176; 12'd173: toneL = 32'd1176; 
                12'd174: toneL = 32'd1176; 12'd175: toneL = `sil; 
                12'd176: toneL = 32'd1048; 12'd177: toneL = 32'd1048; 
                12'd178: toneL = 32'd1048; 12'd179: toneL = `sil; 
                12'd180: toneL = 32'd880; 12'd181: toneL = 32'd880; 
                12'd182: toneL = 32'd880; 12'd183: toneL = `sil; 
                12'd184: toneL = 32'd698; 12'd185: toneL = 32'd698; 
                12'd186: toneL = 32'd698; 12'd187: toneL = `sil; 
                12'd188: toneL = 32'd588; 12'd189: toneL = 32'd588; 
                12'd190: toneL = 32'd588; 12'd191: toneL = `sil; 
                12'd192: toneL = 32'd466; 12'd193: toneL = 32'd466; 
                12'd194: toneL = 32'd466; 12'd195: toneL = `sil; 
                12'd196: toneL = 32'd588; 12'd197: toneL = 32'd588; 
                12'd198: toneL = 32'd588; 12'd199: toneL = `sil; 
                12'd200: toneL = 32'd698; 12'd201: toneL = 32'd698; 
                12'd202: toneL = 32'd698; 12'd203: toneL = `sil; 
                12'd204: toneL = 32'd932; 12'd205: toneL = 32'd932; 
                12'd206: toneL = 32'd932; 12'd207: toneL = `sil; 
                12'd208: toneL = 32'd1176; 12'd209: toneL = 32'd1176; 
                12'd210: toneL = 32'd1176; 12'd211: toneL = `sil; 
                12'd212: toneL = 32'd1396; 12'd213: toneL = 32'd1396; 
                12'd214: toneL = 32'd1396; 12'd215: toneL = `sil; 
                12'd216: toneL = 32'd1864; 12'd217: toneL = 32'd1864; 
                12'd218: toneL = 32'd1864; 12'd219: toneL = `sil; 
                12'd220: toneL = 32'd2096; 12'd221: toneL = 32'd2096; 
                12'd222: toneL = 32'd2096; 12'd223: toneL = `sil; 
                12'd224: toneL = 32'd2096; 12'd225: toneL = 32'd2096; 
                12'd226: toneL = 32'd2096; 12'd227: toneL = `sil; 
                12'd228: toneL = 32'd1864; 12'd229: toneL = 32'd1864; 
                12'd230: toneL = 32'd1864; 12'd231: toneL = `sil; 
                12'd232: toneL = 32'd1396; 12'd233: toneL = 32'd1396; 
                12'd234: toneL = 32'd1396; 12'd235: toneL = `sil; 
                12'd236: toneL = 32'd1176; 12'd237: toneL = 32'd1176; 
                12'd238: toneL = 32'd1176; 12'd239: toneL = `sil; 
                12'd240: toneL = 32'd1048; 12'd241: toneL = 32'd1048; 
                12'd242: toneL = 32'd1048; 12'd243: toneL = `sil; 
                12'd244: toneL = 32'd932; 12'd245: toneL = 32'd932; 
                12'd246: toneL = 32'd932; 12'd247: toneL = `sil; 
                12'd248: toneL = 32'd698; 12'd249: toneL = 32'd698; 
                12'd250: toneL = 32'd698; 12'd251: toneL = `sil; 
                12'd252: toneL = 32'd588; 12'd253: toneL = 32'd588; 
                12'd254: toneL = 32'd588; 12'd255: toneL = `sil; 
                12'd256: toneL = 32'd524; 12'd257: toneL = 32'd524; 
                12'd258: toneL = 32'd524; 12'd259: toneL = `sil; 
                12'd260: toneL = 32'd698; 12'd261: toneL = 32'd698; 
                12'd262: toneL = 32'd698; 12'd263: toneL = `sil; 
                12'd264: toneL = 32'd880; 12'd265: toneL = 32'd880; 
                12'd266: toneL = 32'd880; 12'd267: toneL = `sil; 
                12'd268: toneL = 32'd1048; 12'd269: toneL = 32'd1048; 
                12'd270: toneL = 32'd1048; 12'd271: toneL = `sil; 
                12'd272: toneL = 32'd1048; 12'd273: toneL = 32'd1048; 
                12'd274: toneL = 32'd1048; 12'd275: toneL = `sil; 
                12'd276: toneL = 32'd1396; 12'd277: toneL = 32'd1396; 
                12'd278: toneL = 32'd1396; 12'd279: toneL = `sil; 
                12'd280: toneL = 32'd1760; 12'd281: toneL = 32'd1760; 
                12'd282: toneL = 32'd1760; 12'd283: toneL = `sil; 
                12'd284: toneL = 32'd2096; 12'd285: toneL = 32'd2096; 
                12'd286: toneL = 32'd2096; 12'd287: toneL = `sil; 
                12'd288: toneL = 32'd2096; 12'd289: toneL = 32'd2096; 
                12'd290: toneL = 32'd2096; 12'd291: toneL = `sil; 
                12'd292: toneL = 32'd1760; 12'd293: toneL = 32'd1760; 
                12'd294: toneL = 32'd1760; 12'd295: toneL = `sil; 
                12'd296: toneL = 32'd1396; 12'd297: toneL = 32'd1396; 
                12'd298: toneL = 32'd1396; 12'd299: toneL = `sil; 
                12'd300: toneL = 32'd1048; 12'd301: toneL = 32'd1048; 
                12'd302: toneL = 32'd1048; 12'd303: toneL = `sil; 
                12'd304: toneL = 32'd1048; 12'd305: toneL = 32'd1048; 
                12'd306: toneL = 32'd1048; 12'd307: toneL = `sil; 
                12'd308: toneL = 32'd880; 12'd309: toneL = 32'd880; 
                12'd310: toneL = 32'd880; 12'd311: toneL = `sil; 
                12'd312: toneL = 32'd698; 12'd313: toneL = 32'd698; 
                12'd314: toneL = 32'd698; 12'd315: toneL = `sil; 
                12'd316: toneL = 32'd524; 12'd317: toneL = 32'd524; 
                12'd318: toneL = 32'd524; 12'd319: toneL = `sil; 
                12'd320: toneL = 32'd524; 12'd321: toneL = 32'd524; 
                12'd322: toneL = 32'd524; 12'd323: toneL = `sil; 
                12'd324: toneL = 32'd660; 12'd325: toneL = 32'd660; 
                12'd326: toneL = 32'd660; 12'd327: toneL = `sil; 
                12'd328: toneL = 32'd784; 12'd329: toneL = 32'd784; 
                12'd330: toneL = 32'd784; 12'd331: toneL = `sil; 
                12'd332: toneL = 32'd1048; 12'd333: toneL = 32'd1048; 
                12'd334: toneL = 32'd1048; 12'd335: toneL = `sil; 
                12'd336: toneL = 32'd1048; 12'd337: toneL = 32'd1048; 
                12'd338: toneL = 32'd1048; 12'd339: toneL = `sil; 
                12'd340: toneL = 32'd1320; 12'd341: toneL = 32'd1320; 
                12'd342: toneL = 32'd1320; 12'd343: toneL = `sil; 
                12'd344: toneL = 32'd1568; 12'd345: toneL = 32'd1568; 
                12'd346: toneL = 32'd1568; 12'd347: toneL = `sil; 
                12'd348: toneL = 32'd2096; 12'd349: toneL = 32'd2096; 
                12'd350: toneL = 32'd2096; 12'd351: toneL = `sil; 
                12'd352: toneL = 32'd2096; 12'd353: toneL = 32'd2096; 
                12'd354: toneL = 32'd2096; 12'd355: toneL = `sil; 
                12'd356: toneL = 32'd1568; 12'd357: toneL = 32'd1568; 
                12'd358: toneL = 32'd1568; 12'd359: toneL = `sil; 
                12'd360: toneL = 32'd1320; 12'd361: toneL = 32'd1320; 
                12'd362: toneL = 32'd1320; 12'd363: toneL = `sil; 
                12'd364: toneL = 32'd1048; 12'd365: toneL = 32'd1048; 
                12'd366: toneL = 32'd1048; 12'd367: toneL = `sil; 
                12'd368: toneL = 32'd1048; 12'd369: toneL = 32'd1048; 
                12'd370: toneL = 32'd1048; 12'd371: toneL = `sil; 
                12'd372: toneL = 32'd784; 12'd373: toneL = 32'd784; 
                12'd374: toneL = 32'd784; 12'd375: toneL = `sil; 
                12'd376: toneL = 32'd660; 12'd377: toneL = 32'd660; 
                12'd378: toneL = 32'd660; 12'd379: toneL = `sil; 
                12'd380: toneL = 32'd524; 12'd381: toneL = 32'd524; 
                12'd382: toneL = 32'd524; 12'd383: toneL = `sil; 
                12'd384: toneL = 32'd588; 12'd385: toneL = 32'd588; 
                12'd386: toneL = 32'd588; 12'd387: toneL = `sil; 
                12'd388: toneL = 32'd698; 12'd389: toneL = 32'd698; 
                12'd390: toneL = 32'd698; 12'd391: toneL = `sil; 
                12'd392: toneL = 32'd880; 12'd393: toneL = 32'd880; 
                12'd394: toneL = 32'd880; 12'd395: toneL = `sil; 
                12'd396: toneL = 32'd1048; 12'd397: toneL = 32'd1048; 
                12'd398: toneL = 32'd1048; 12'd399: toneL = `sil; 
                12'd400: toneL = 32'd1176; 12'd401: toneL = 32'd1176; 
                12'd402: toneL = 32'd1176; 12'd403: toneL = `sil; 
                12'd404: toneL = 32'd1396; 12'd405: toneL = 32'd1396; 
                12'd406: toneL = 32'd1396; 12'd407: toneL = `sil; 
                12'd408: toneL = 32'd1760; 12'd409: toneL = 32'd1760; 
                12'd410: toneL = 32'd1760; 12'd411: toneL = `sil; 
                12'd412: toneL = 32'd2096; 12'd413: toneL = 32'd2096; 
                12'd414: toneL = 32'd2096; 12'd415: toneL = `sil; 
                12'd416: toneL = 32'd2096; 12'd417: toneL = 32'd2096; 
                12'd418: toneL = 32'd2096; 12'd419: toneL = `sil; 
                12'd420: toneL = 32'd1760; 12'd421: toneL = 32'd1760; 
                12'd422: toneL = 32'd1760; 12'd423: toneL = `sil; 
                12'd424: toneL = 32'd1396; 12'd425: toneL = 32'd1396; 
                12'd426: toneL = 32'd1396; 12'd427: toneL = `sil; 
                12'd428: toneL = 32'd1176; 12'd429: toneL = 32'd1176; 
                12'd430: toneL = 32'd1176; 12'd431: toneL = `sil; 
                12'd432: toneL = 32'd1048; 12'd433: toneL = 32'd1048; 
                12'd434: toneL = 32'd1048; 12'd435: toneL = `sil; 
                12'd436: toneL = 32'd880; 12'd437: toneL = 32'd880; 
                12'd438: toneL = 32'd880; 12'd439: toneL = `sil; 
                12'd440: toneL = 32'd698; 12'd441: toneL = 32'd698; 
                12'd442: toneL = 32'd698; 12'd443: toneL = `sil; 
                12'd444: toneL = 32'd588; 12'd445: toneL = 32'd588; 
                12'd446: toneL = 32'd588; 12'd447: toneL = `sil; 
                12'd448: toneL = 32'd466; 12'd449: toneL = 32'd466; 
                12'd450: toneL = 32'd466; 12'd451: toneL = `sil; 
                12'd452: toneL = 32'd588; 12'd453: toneL = 32'd588; 
                12'd454: toneL = 32'd588; 12'd455: toneL = `sil; 
                12'd456: toneL = 32'd698; 12'd457: toneL = 32'd698; 
                12'd458: toneL = 32'd698; 12'd459: toneL = `sil; 
                12'd460: toneL = 32'd932; 12'd461: toneL = 32'd932; 
                12'd462: toneL = 32'd932; 12'd463: toneL = `sil; 
                12'd464: toneL = 32'd1176; 12'd465: toneL = 32'd1176; 
                12'd466: toneL = 32'd1176; 12'd467: toneL = `sil; 
                12'd468: toneL = 32'd1396; 12'd469: toneL = 32'd1396; 
                12'd470: toneL = 32'd1396; 12'd471: toneL = `sil; 
                12'd472: toneL = 32'd1864; 12'd473: toneL = 32'd1864; 
                12'd474: toneL = 32'd1864; 12'd475: toneL = `sil; 
                12'd476: toneL = 32'd2096; 12'd477: toneL = 32'd2096; 
                12'd478: toneL = 32'd2096; 12'd479: toneL = `sil; 
                12'd480: toneL = 32'd2096; 12'd481: toneL = 32'd2096; 
                12'd482: toneL = 32'd2096; 12'd483: toneL = `sil; 
                12'd484: toneL = 32'd1864; 12'd485: toneL = 32'd1864; 
                12'd486: toneL = 32'd1864; 12'd487: toneL = `sil; 
                12'd488: toneL = 32'd1396; 12'd489: toneL = 32'd1396; 
                12'd490: toneL = 32'd1396; 12'd491: toneL = `sil; 
                12'd492: toneL = 32'd1176; 12'd493: toneL = 32'd1176; 
                12'd494: toneL = 32'd1176; 12'd495: toneL = `sil; 
                12'd496: toneL = 32'd1048; 12'd497: toneL = 32'd1048; 
                12'd498: toneL = 32'd1048; 12'd499: toneL = `sil; 
                12'd500: toneL = 32'd932; 12'd501: toneL = 32'd932; 
                12'd502: toneL = 32'd932; 12'd503: toneL = `sil; 
                12'd504: toneL = 32'd698; 12'd505: toneL = 32'd698; 
                12'd506: toneL = 32'd698; 12'd507: toneL = `sil; 
                12'd508: toneL = 32'd588; 12'd509: toneL = 32'd588; 
                12'd510: toneL = 32'd588; 12'd511: toneL = `sil; 
                12'd512: toneL = 32'd524; 12'd513: toneL = 32'd524; 
                12'd514: toneL = 32'd524; 12'd515: toneL = `sil; 
                12'd516: toneL = 32'd698; 12'd517: toneL = 32'd698; 
                12'd518: toneL = 32'd698; 12'd519: toneL = `sil; 
                12'd520: toneL = 32'd880; 12'd521: toneL = 32'd880; 
                12'd522: toneL = 32'd880; 12'd523: toneL = `sil; 
                12'd524: toneL = 32'd1048; 12'd525: toneL = 32'd1048; 
                12'd526: toneL = 32'd1048; 12'd527: toneL = `sil; 
                12'd528: toneL = 32'd1048; 12'd529: toneL = 32'd1048; 
                12'd530: toneL = 32'd1048; 12'd531: toneL = `sil; 
                12'd532: toneL = 32'd1396; 12'd533: toneL = 32'd1396; 
                12'd534: toneL = 32'd1396; 12'd535: toneL = `sil; 
                12'd536: toneL = 32'd1760; 12'd537: toneL = 32'd1760; 
                12'd538: toneL = 32'd1760; 12'd539: toneL = `sil; 
                12'd540: toneL = 32'd2096; 12'd541: toneL = 32'd2096; 
                12'd542: toneL = 32'd2096; 12'd543: toneL = `sil; 
                12'd544: toneL = 32'd2096; 12'd545: toneL = 32'd2096; 
                12'd546: toneL = 32'd2096; 12'd547: toneL = `sil; 
                12'd548: toneL = 32'd1760; 12'd549: toneL = 32'd1760; 
                12'd550: toneL = 32'd1760; 12'd551: toneL = `sil; 
                12'd552: toneL = 32'd1396; 12'd553: toneL = 32'd1396; 
                12'd554: toneL = 32'd1396; 12'd555: toneL = `sil; 
                12'd556: toneL = 32'd1048; 12'd557: toneL = 32'd1048; 
                12'd558: toneL = 32'd1048; 12'd559: toneL = `sil; 
                12'd560: toneL = 32'd1048; 12'd561: toneL = 32'd1048; 
                12'd562: toneL = 32'd1048; 12'd563: toneL = `sil; 
                12'd564: toneL = 32'd880; 12'd565: toneL = 32'd880; 
                12'd566: toneL = 32'd880; 12'd567: toneL = `sil; 
                12'd568: toneL = 32'd698; 12'd569: toneL = 32'd698; 
                12'd570: toneL = 32'd698; 12'd571: toneL = `sil; 
                12'd572: toneL = 32'd524; 12'd573: toneL = 32'd524; 
                12'd574: toneL = 32'd524; 12'd575: toneL = `sil; 
                12'd576: toneL = 32'd524; 12'd577: toneL = 32'd524; 
                12'd578: toneL = 32'd524; 12'd579: toneL = `sil; 
                12'd580: toneL = 32'd660; 12'd581: toneL = 32'd660; 
                12'd582: toneL = 32'd660; 12'd583: toneL = `sil; 
                12'd584: toneL = 32'd784; 12'd585: toneL = 32'd784; 
                12'd586: toneL = 32'd784; 12'd587: toneL = `sil; 
                12'd588: toneL = 32'd1048; 12'd589: toneL = 32'd1048; 
                12'd590: toneL = 32'd1048; 12'd591: toneL = `sil; 
                12'd592: toneL = 32'd1048; 12'd593: toneL = 32'd1048; 
                12'd594: toneL = 32'd1048; 12'd595: toneL = `sil; 
                12'd596: toneL = 32'd1320; 12'd597: toneL = 32'd1320; 
                12'd598: toneL = 32'd1320; 12'd599: toneL = `sil; 
                12'd600: toneL = 32'd1568; 12'd601: toneL = 32'd1568; 
                12'd602: toneL = 32'd1568; 12'd603: toneL = `sil; 
                12'd604: toneL = 32'd2096; 12'd605: toneL = 32'd2096; 
                12'd606: toneL = 32'd2096; 12'd607: toneL = `sil; 
                12'd608: toneL = 32'd2096; 12'd609: toneL = 32'd2096; 
                12'd610: toneL = 32'd2096; 12'd611: toneL = `sil; 
                12'd612: toneL = 32'd1568; 12'd613: toneL = 32'd1568; 
                12'd614: toneL = 32'd1568; 12'd615: toneL = `sil; 
                12'd616: toneL = 32'd1320; 12'd617: toneL = 32'd1320; 
                12'd618: toneL = 32'd1320; 12'd619: toneL = `sil; 
                12'd620: toneL = 32'd1048; 12'd621: toneL = 32'd1048; 
                12'd622: toneL = 32'd1048; 12'd623: toneL = `sil; 
                12'd624: toneL = 32'd1048; 12'd625: toneL = 32'd1048; 
                12'd626: toneL = 32'd1048; 12'd627: toneL = `sil; 
                12'd628: toneL = 32'd784; 12'd629: toneL = 32'd784; 
                12'd630: toneL = 32'd784; 12'd631: toneL = `sil; 
                12'd632: toneL = 32'd660; 12'd633: toneL = 32'd660; 
                12'd634: toneL = 32'd660; 12'd635: toneL = `sil; 
                12'd636: toneL = 32'd524; 12'd637: toneL = 32'd524; 
                12'd638: toneL = 32'd524; 12'd639: toneL = `sil; 
                12'd640: toneL = 32'd588; 12'd641: toneL = 32'd588; 
                12'd642: toneL = 32'd588; 12'd643: toneL = `sil; 
                12'd644: toneL = 32'd698; 12'd645: toneL = 32'd698; 
                12'd646: toneL = 32'd698; 12'd647: toneL = `sil; 
                12'd648: toneL = 32'd880; 12'd649: toneL = 32'd880; 
                12'd650: toneL = 32'd880; 12'd651: toneL = `sil; 
                12'd652: toneL = 32'd1048; 12'd653: toneL = 32'd1048; 
                12'd654: toneL = 32'd1048; 12'd655: toneL = `sil; 
                12'd656: toneL = 32'd1176; 12'd657: toneL = 32'd1176; 
                12'd658: toneL = 32'd1176; 12'd659: toneL = `sil; 
                12'd660: toneL = 32'd1396; 12'd661: toneL = 32'd1396; 
                12'd662: toneL = 32'd1396; 12'd663: toneL = `sil; 
                12'd664: toneL = 32'd1760; 12'd665: toneL = 32'd1760; 
                12'd666: toneL = 32'd1760; 12'd667: toneL = `sil; 
                12'd668: toneL = 32'd2096; 12'd669: toneL = 32'd2096; 
                12'd670: toneL = 32'd2096; 12'd671: toneL = `sil; 
                12'd672: toneL = 32'd2096; 12'd673: toneL = 32'd2096; 
                12'd674: toneL = 32'd2096; 12'd675: toneL = `sil; 
                12'd676: toneL = 32'd1760; 12'd677: toneL = 32'd1760; 
                12'd678: toneL = 32'd1760; 12'd679: toneL = `sil; 
                12'd680: toneL = 32'd1396; 12'd681: toneL = 32'd1396; 
                12'd682: toneL = 32'd1396; 12'd683: toneL = `sil; 
                12'd684: toneL = 32'd1176; 12'd685: toneL = 32'd1176; 
                12'd686: toneL = 32'd1176; 12'd687: toneL = `sil; 
                12'd688: toneL = 32'd1048; 12'd689: toneL = 32'd1048; 
                12'd690: toneL = 32'd1048; 12'd691: toneL = `sil; 
                12'd692: toneL = 32'd880; 12'd693: toneL = 32'd880; 
                12'd694: toneL = 32'd880; 12'd695: toneL = `sil; 
                12'd696: toneL = 32'd698; 12'd697: toneL = 32'd698; 
                12'd698: toneL = 32'd698; 12'd699: toneL = `sil; 
                12'd700: toneL = 32'd588; 12'd701: toneL = 32'd588; 
                12'd702: toneL = 32'd588; 12'd703: toneL = `sil; 
                12'd704: toneL = 32'd466; 12'd705: toneL = 32'd466; 
                12'd706: toneL = 32'd466; 12'd707: toneL = `sil; 
                12'd708: toneL = 32'd588; 12'd709: toneL = 32'd588; 
                12'd710: toneL = 32'd588; 12'd711: toneL = `sil; 
                12'd712: toneL = 32'd698; 12'd713: toneL = 32'd698; 
                12'd714: toneL = 32'd698; 12'd715: toneL = `sil; 
                12'd716: toneL = 32'd932; 12'd717: toneL = 32'd932; 
                12'd718: toneL = 32'd932; 12'd719: toneL = `sil; 
                12'd720: toneL = 32'd1176; 12'd721: toneL = 32'd1176; 
                12'd722: toneL = 32'd1176; 12'd723: toneL = `sil; 
                12'd724: toneL = 32'd1396; 12'd725: toneL = 32'd1396; 
                12'd726: toneL = 32'd1396; 12'd727: toneL = `sil; 
                12'd728: toneL = 32'd1864; 12'd729: toneL = 32'd1864; 
                12'd730: toneL = 32'd1864; 12'd731: toneL = `sil; 
                12'd732: toneL = 32'd2096; 12'd733: toneL = 32'd2096; 
                12'd734: toneL = 32'd2096; 12'd735: toneL = `sil; 
                12'd736: toneL = 32'd2096; 12'd737: toneL = 32'd2096; 
                12'd738: toneL = 32'd2096; 12'd739: toneL = `sil; 
                12'd740: toneL = 32'd1864; 12'd741: toneL = 32'd1864; 
                12'd742: toneL = 32'd1864; 12'd743: toneL = `sil; 
                12'd744: toneL = 32'd1396; 12'd745: toneL = 32'd1396; 
                12'd746: toneL = 32'd1396; 12'd747: toneL = `sil; 
                12'd748: toneL = 32'd1176; 12'd749: toneL = 32'd1176; 
                12'd750: toneL = 32'd1176; 12'd751: toneL = `sil; 
                12'd752: toneL = 32'd1048; 12'd753: toneL = 32'd1048; 
                12'd754: toneL = 32'd1048; 12'd755: toneL = `sil; 
                12'd756: toneL = 32'd932; 12'd757: toneL = 32'd932; 
                12'd758: toneL = 32'd932; 12'd759: toneL = `sil; 
                12'd760: toneL = 32'd698; 12'd761: toneL = 32'd698; 
                12'd762: toneL = 32'd698; 12'd763: toneL = `sil; 
                12'd764: toneL = 32'd588; 12'd765: toneL = 32'd588; 
                12'd766: toneL = 32'd588; 12'd767: toneL = `sil; 
                12'd768: toneL = 32'd524; 12'd769: toneL = 32'd524; 
                12'd770: toneL = 32'd524; 12'd771: toneL = `sil; 
                12'd772: toneL = 32'd698; 12'd773: toneL = 32'd698; 
                12'd774: toneL = 32'd698; 12'd775: toneL = `sil; 
                12'd776: toneL = 32'd880; 12'd777: toneL = 32'd880; 
                12'd778: toneL = 32'd880; 12'd779: toneL = `sil; 
                12'd780: toneL = 32'd1048; 12'd781: toneL = 32'd1048; 
                12'd782: toneL = 32'd1048; 12'd783: toneL = `sil; 
                12'd784: toneL = 32'd1048; 12'd785: toneL = 32'd1048; 
                12'd786: toneL = 32'd1048; 12'd787: toneL = `sil; 
                12'd788: toneL = 32'd1396; 12'd789: toneL = 32'd1396; 
                12'd790: toneL = 32'd1396; 12'd791: toneL = `sil; 
                12'd792: toneL = 32'd1760; 12'd793: toneL = 32'd1760; 
                12'd794: toneL = 32'd1760; 12'd795: toneL = `sil; 
                12'd796: toneL = 32'd2096; 12'd797: toneL = 32'd2096; 
                12'd798: toneL = 32'd2096; 12'd799: toneL = `sil; 
                12'd800: toneL = 32'd2096; 12'd801: toneL = 32'd2096; 
                12'd802: toneL = 32'd2096; 12'd803: toneL = `sil; 
                12'd804: toneL = 32'd1760; 12'd805: toneL = 32'd1760; 
                12'd806: toneL = 32'd1760; 12'd807: toneL = `sil; 
                12'd808: toneL = 32'd1396; 12'd809: toneL = 32'd1396; 
                12'd810: toneL = 32'd1396; 12'd811: toneL = `sil; 
                12'd812: toneL = 32'd1048; 12'd813: toneL = 32'd1048; 
                12'd814: toneL = 32'd1048; 12'd815: toneL = `sil; 
                12'd816: toneL = 32'd1048; 12'd817: toneL = 32'd1048; 
                12'd818: toneL = 32'd1048; 12'd819: toneL = `sil; 
                12'd820: toneL = 32'd880; 12'd821: toneL = 32'd880; 
                12'd822: toneL = 32'd880; 12'd823: toneL = `sil; 
                12'd824: toneL = 32'd698; 12'd825: toneL = 32'd698; 
                12'd826: toneL = 32'd698; 12'd827: toneL = `sil; 
                12'd828: toneL = 32'd524; 12'd829: toneL = 32'd524; 
                12'd830: toneL = 32'd524; 12'd831: toneL = `sil; 
                12'd832: toneL = 32'd524; 12'd833: toneL = 32'd524; 
                12'd834: toneL = 32'd524; 12'd835: toneL = `sil; 
                12'd836: toneL = 32'd660; 12'd837: toneL = 32'd660; 
                12'd838: toneL = 32'd660; 12'd839: toneL = `sil; 
                12'd840: toneL = 32'd784; 12'd841: toneL = 32'd784; 
                12'd842: toneL = 32'd784; 12'd843: toneL = `sil; 
                12'd844: toneL = 32'd1048; 12'd845: toneL = 32'd1048; 
                12'd846: toneL = 32'd1048; 12'd847: toneL = `sil; 
                12'd848: toneL = 32'd1048; 12'd849: toneL = 32'd1048; 
                12'd850: toneL = 32'd1048; 12'd851: toneL = `sil; 
                12'd852: toneL = 32'd1320; 12'd853: toneL = 32'd1320; 
                12'd854: toneL = 32'd1320; 12'd855: toneL = `sil; 
                12'd856: toneL = 32'd1568; 12'd857: toneL = 32'd1568; 
                12'd858: toneL = 32'd1568; 12'd859: toneL = `sil; 
                12'd860: toneL = 32'd2096; 12'd861: toneL = 32'd2096; 
                12'd862: toneL = 32'd2096; 12'd863: toneL = `sil; 
                12'd864: toneL = 32'd2096; 12'd865: toneL = 32'd2096; 
                12'd866: toneL = 32'd2096; 12'd867: toneL = `sil; 
                12'd868: toneL = 32'd1568; 12'd869: toneL = 32'd1568; 
                12'd870: toneL = 32'd1568; 12'd871: toneL = `sil; 
                12'd872: toneL = 32'd1320; 12'd873: toneL = 32'd1320; 
                12'd874: toneL = 32'd1320; 12'd875: toneL = `sil; 
                12'd876: toneL = 32'd1048; 12'd877: toneL = 32'd1048; 
                12'd878: toneL = 32'd1048; 12'd879: toneL = `sil; 
                12'd880: toneL = 32'd1048; 12'd881: toneL = 32'd1048; 
                12'd882: toneL = 32'd1048; 12'd883: toneL = `sil; 
                12'd884: toneL = 32'd784; 12'd885: toneL = 32'd784; 
                12'd886: toneL = 32'd784; 12'd887: toneL = `sil; 
                12'd888: toneL = 32'd660; 12'd889: toneL = 32'd660; 
                12'd890: toneL = 32'd660; 12'd891: toneL = `sil; 
                12'd892: toneL = 32'd524; 12'd893: toneL = 32'd524; 
                12'd894: toneL = 32'd524; 12'd895: toneL = `sil; 
                12'd896: toneL = 32'd588; 12'd897: toneL = 32'd588; 
                12'd898: toneL = 32'd588; 12'd899: toneL = `sil; 
                12'd900: toneL = 32'd698; 12'd901: toneL = 32'd698; 
                12'd902: toneL = 32'd698; 12'd903: toneL = `sil; 
                12'd904: toneL = 32'd880; 12'd905: toneL = 32'd880; 
                12'd906: toneL = 32'd880; 12'd907: toneL = `sil; 
                12'd908: toneL = 32'd1048; 12'd909: toneL = 32'd1048; 
                12'd910: toneL = 32'd1048; 12'd911: toneL = `sil; 
                12'd912: toneL = 32'd1176; 12'd913: toneL = 32'd1176; 
                12'd914: toneL = 32'd1176; 12'd915: toneL = `sil; 
                12'd916: toneL = 32'd1396; 12'd917: toneL = 32'd1396; 
                12'd918: toneL = 32'd1396; 12'd919: toneL = `sil; 
                12'd920: toneL = 32'd1760; 12'd921: toneL = 32'd1760; 
                12'd922: toneL = 32'd1760; 12'd923: toneL = `sil; 
                12'd924: toneL = 32'd2096; 12'd925: toneL = 32'd2096; 
                12'd926: toneL = 32'd2096; 12'd927: toneL = `sil; 
                12'd928: toneL = 32'd2096; 12'd929: toneL = 32'd2096; 
                12'd930: toneL = 32'd2096; 12'd931: toneL = `sil; 
                12'd932: toneL = 32'd1760; 12'd933: toneL = 32'd1760; 
                12'd934: toneL = 32'd1760; 12'd935: toneL = `sil; 
                12'd936: toneL = 32'd1396; 12'd937: toneL = 32'd1396; 
                12'd938: toneL = 32'd1396; 12'd939: toneL = `sil; 
                12'd940: toneL = 32'd1176; 12'd941: toneL = 32'd1176; 
                12'd942: toneL = 32'd1176; 12'd943: toneL = `sil; 
                12'd944: toneL = 32'd1048; 12'd945: toneL = 32'd1048; 
                12'd946: toneL = 32'd1048; 12'd947: toneL = `sil; 
                12'd948: toneL = 32'd880; 12'd949: toneL = 32'd880; 
                12'd950: toneL = 32'd880; 12'd951: toneL = `sil; 
                12'd952: toneL = 32'd698; 12'd953: toneL = 32'd698; 
                12'd954: toneL = 32'd698; 12'd955: toneL = `sil; 
                12'd956: toneL = 32'd588; 12'd957: toneL = 32'd588; 
                12'd958: toneL = 32'd588; 12'd959: toneL = `sil; 
                12'd960: toneL = 32'd466; 12'd961: toneL = 32'd466; 
                12'd962: toneL = 32'd466; 12'd963: toneL = `sil; 
                12'd964: toneL = 32'd588; 12'd965: toneL = 32'd588; 
                12'd966: toneL = 32'd588; 12'd967: toneL = `sil; 
                12'd968: toneL = 32'd698; 12'd969: toneL = 32'd698; 
                12'd970: toneL = 32'd698; 12'd971: toneL = `sil; 
                12'd972: toneL = 32'd932; 12'd973: toneL = 32'd932; 
                12'd974: toneL = 32'd932; 12'd975: toneL = `sil; 
                12'd976: toneL = 32'd1176; 12'd977: toneL = 32'd1176; 
                12'd978: toneL = 32'd1176; 12'd979: toneL = `sil; 
                12'd980: toneL = 32'd1396; 12'd981: toneL = 32'd1396; 
                12'd982: toneL = 32'd1396; 12'd983: toneL = `sil; 
                12'd984: toneL = 32'd1864; 12'd985: toneL = 32'd1864; 
                12'd986: toneL = 32'd1864; 12'd987: toneL = `sil; 
                12'd988: toneL = 32'd2096; 12'd989: toneL = 32'd2096; 
                12'd990: toneL = 32'd2096; 12'd991: toneL = `sil; 
                12'd992: toneL = 32'd2096; 12'd993: toneL = 32'd2096; 
                12'd994: toneL = 32'd2096; 12'd995: toneL = `sil; 
                12'd996: toneL = 32'd1864; 12'd997: toneL = 32'd1864; 
                12'd998: toneL = 32'd1864; 12'd999: toneL = `sil; 
                12'd1000: toneL = 32'd1396; 12'd1001: toneL = 32'd1396; 
                12'd1002: toneL = 32'd1396; 12'd1003: toneL = `sil; 
                12'd1004: toneL = 32'd1176; 12'd1005: toneL = 32'd1176; 
                12'd1006: toneL = 32'd1176; 12'd1007: toneL = `sil; 
                12'd1008: toneL = 32'd1048; 12'd1009: toneL = 32'd1048; 
                12'd1010: toneL = 32'd1048; 12'd1011: toneL = `sil; 
                12'd1012: toneL = 32'd932; 12'd1013: toneL = 32'd932; 
                12'd1014: toneL = 32'd932; 12'd1015: toneL = `sil; 
                12'd1016: toneL = 32'd698; 12'd1017: toneL = 32'd698; 
                12'd1018: toneL = 32'd698; 12'd1019: toneL = `sil; 
                12'd1020: toneL = 32'd588; 12'd1021: toneL = 32'd588; 
                12'd1022: toneL = 32'd588; 12'd1023: toneL = `sil; 



                default : toneL = `sil;
            endcase
        end
        else /*if (state_for_L_ch == 1'b1*//*waiting_playing*//*)*/ begin
            case(ibeatNum)
                12'd0: toneL = 32'd392; 12'd1: toneL = 32'd392; 
                12'd2: toneL = 32'd392; 12'd3: toneL = 32'd392; 
                12'd4: toneL = 32'd392; 12'd5: toneL = 32'd392;
                12'd6: toneL = 32'd415; 12'd7: toneL = 32'd415;
                12'd8: toneL = 32'd440; 12'd9: toneL = 32'd440; 
                12'd10: toneL = 32'd440; 12'd11: toneL = 32'd440; 
                12'd12: toneL = 32'd440; 12'd13: toneL = 32'd440; 
                12'd14: toneL = 32'd440; 12'd15: toneL = 32'd440; 
                12'd16: toneL = 32'd440; 12'd17: toneL = 32'd440; 
                12'd18: toneL = 32'd440; 12'd19: toneL = 32'd440; 
                12'd20: toneL = 32'd440; 12'd21: toneL = 32'd440; 
                12'd22: toneL = 32'd440; 12'd23: toneL = 32'd440; 
                12'd24: toneL = 32'd440; 12'd25: toneL = 32'd440; 
                12'd26: toneL = 32'd440; 12'd27: toneL = 32'd440; 
                12'd28: toneL = 32'd440; 12'd29: toneL = 32'd440; 
                12'd30: toneL = 32'd440; 12'd31: toneL = 32'd440; 
                12'd32: toneL = 32'd440; 12'd33: toneL = 32'd440; 
                12'd34: toneL = 32'd440; 12'd35: toneL = 32'd440; 
                12'd36: toneL = 32'd440; 12'd37: toneL = 32'd440; 
                12'd38: toneL = 32'd440; 12'd39: toneL = 32'd440; 
                12'd40: toneL = 32'd440; 12'd41: toneL = 32'd440; 
                12'd42: toneL = 32'd440; 12'd43: toneL = 32'd440; 
                12'd44: toneL = 32'd440; 12'd45: toneL = 32'd440; 
                12'd46: toneL = 32'd392; 12'd47: toneL = 32'd392;
                12'd48: toneL = 32'd440; 12'd49: toneL = 32'd440; 
                12'd50: toneL = 32'd440; 12'd51: toneL = 32'd440; 
                12'd52: toneL = 32'd440; 12'd53: toneL = 32'd440;
                12'd54: toneL = 32'd392; 12'd55: toneL = 32'd392;
                12'd56: toneL = 32'd440; 12'd57: toneL = 32'd440; 
                12'd58: toneL = 32'd440; 12'd59: toneL = 32'd440; 
                12'd60: toneL = 32'd440; 12'd61: toneL = 32'd440; 
                12'd62: toneL = 32'd392; 12'd63: toneL = 32'd392;
                12'd64: toneL = 32'd330; 12'd65: toneL = 32'd330; 
                12'd66: toneL = 32'd330; 12'd67: toneL = 32'd330; 
                12'd68: toneL = 32'd330; 12'd69: toneL = 32'd330; 
                12'd70: toneL = 32'd262; 12'd71: toneL = 32'd262;
                12'd72: toneL = 32'd440; 12'd73: toneL = 32'd440; 
                12'd74: toneL = 32'd440; 12'd75: toneL = 32'd440; 
                12'd76: toneL = 32'd440; 12'd77: toneL = 32'd440; 
                12'd78: toneL = 32'd440; 12'd79: toneL = 32'd440; 
                12'd80: toneL = 32'd440; 12'd81: toneL = 32'd440; 
                12'd82: toneL = 32'd440; 12'd83: toneL = 32'd440; 
                12'd84: toneL = 32'd440; 12'd85: toneL = 32'd440; 
                12'd86: toneL = 32'd440; 12'd87: toneL = 32'd440; 
                12'd88: toneL = 32'd440; 12'd89: toneL = 32'd440; 
                12'd90: toneL = 32'd440; 12'd91: toneL = 32'd440; 
                12'd92: toneL = 32'd440; 12'd93: toneL = 32'd440; 
                12'd94: toneL = 32'd440; 12'd95: toneL = 32'd440; 
                12'd96: toneL = 32'd440; 12'd97: toneL = 32'd440; 
                12'd98: toneL = 32'd440; 12'd99: toneL = 32'd440; 
                12'd100: toneL = 32'd440; 12'd101: toneL = 32'd440; 
                12'd102: toneL = 32'd440; 12'd103: toneL = 32'd440; 
                12'd104: toneL = 32'd440; 12'd105: toneL = 32'd440; 
                12'd106: toneL = 32'd440; 12'd107: toneL = 32'd440; 
                12'd108: toneL = 32'd440; 12'd109: toneL = 32'd440; 
                12'd110: toneL = 32'd440; 12'd111: toneL = 32'd440; 
                12'd112: toneL = 32'd440; 12'd113: toneL = 32'd440; 
                12'd114: toneL = 32'd440; 12'd115: toneL = 32'd440; 
                12'd116: toneL = 32'd440; 12'd117: toneL = 32'd440; 
                12'd118: toneL = 32'd440; 12'd119: toneL = 32'd440; 
                12'd120: toneL = 32'd440; 12'd121: toneL = 32'd440; 
                12'd122: toneL = 32'd440; 12'd123: toneL = 32'd440; 
                12'd124: toneL = 32'd440; 12'd125: toneL = 32'd440; 
                12'd126: toneL = 32'd440; 12'd127: toneL = 32'd440; 
                12'd128: toneL = 32'd524; 12'd129: toneL = 32'd524; 
                12'd130: toneL = 32'd524; 12'd131: toneL = 32'd524; 
                12'd132: toneL = 32'd524; 12'd133: toneL = 32'd524;
                12'd134: toneL = 32'd554; 12'd135: toneL = 32'd554;
                12'd136: toneL = 32'd588; 12'd137: toneL = 32'd588; 
                12'd138: toneL = 32'd588; 12'd139: toneL = 32'd588; 
                12'd140: toneL = 32'd588; 12'd141: toneL = 32'd588; 
                12'd142: toneL = 32'd588; 12'd143: toneL = 32'd588; 
                12'd144: toneL = 32'd588; 12'd145: toneL = 32'd588; 
                12'd146: toneL = 32'd588; 12'd147: toneL = 32'd588; 
                12'd148: toneL = 32'd588; 12'd149: toneL = 32'd588; 
                12'd150: toneL = 32'd588; 12'd151: toneL = 32'd588; 
                12'd152: toneL = 32'd588; 12'd153: toneL = 32'd588; 
                12'd154: toneL = 32'd588; 12'd155: toneL = 32'd588; 
                12'd156: toneL = 32'd588; 12'd157: toneL = 32'd588; 
                12'd158: toneL = 32'd588; 12'd159: toneL = 32'd588; 
                12'd160: toneL = 32'd588; 12'd161: toneL = 32'd588; 
                12'd162: toneL = 32'd588; 12'd163: toneL = 32'd588; 
                12'd164: toneL = 32'd588; 12'd165: toneL = 32'd588; 
                12'd166: toneL = 32'd588; 12'd167: toneL = 32'd588; 
                12'd168: toneL = 32'd588; 12'd169: toneL = 32'd588; 
                12'd170: toneL = 32'd588; 12'd171: toneL = 32'd588; 
                12'd172: toneL = 32'd588; 12'd173: toneL = 32'd588; 
                12'd174: toneL = 32'd660; 12'd175: toneL = 32'd660;
                12'd176: toneL = 32'd588; 12'd177: toneL = 32'd588; 
                12'd178: toneL = 32'd588; 12'd179: toneL = 32'd588; 
                12'd180: toneL = 32'd588; 12'd181: toneL = 32'd588; 
                12'd182: toneL = 32'd660; 12'd183: toneL = 32'd660;
                12'd184: toneL = 32'd588; 12'd185: toneL = 32'd588; 
                12'd186: toneL = 32'd588; 12'd187: toneL = 32'd588; 
                12'd188: toneL = 32'd588; 12'd189: toneL = 32'd588; 
                12'd190: toneL = 32'd524; 12'd191: toneL = 32'd524; 
                12'd192: toneL = 32'd524; 12'd193: toneL = 32'd524;
                12'd194: toneL = 32'd415; 12'd195: toneL = 32'd415;
                12'd196: toneL = 32'd349; 12'd197: toneL = 32'd349;
                12'd198: toneL = 32'd588; 12'd199: toneL = 32'd588; 
                12'd200: toneL = 32'd588; 12'd201: toneL = 32'd588; 
                12'd202: toneL = 32'd588; 12'd203: toneL = 32'd588; 
                12'd204: toneL = 32'd588; 12'd205: toneL = 32'd588; 
                12'd206: toneL = 32'd588; 12'd207: toneL = 32'd588; 
                12'd208: toneL = 32'd588; 12'd209: toneL = 32'd588; 
                12'd210: toneL = 32'd588; 12'd211: toneL = 32'd588; 
                12'd212: toneL = 32'd588; 12'd213: toneL = 32'd588; 
                12'd214: toneL = 32'd588; 12'd215: toneL = 32'd588; 
                12'd216: toneL = 32'd588; 12'd217: toneL = 32'd588; 
                12'd218: toneL = 32'd588; 12'd219: toneL = 32'd588; 
                12'd220: toneL = 32'd588; 12'd221: toneL = 32'd588; 
                12'd222: toneL = 32'd588; 12'd223: toneL = 32'd588; 
                12'd224: toneL = 32'd588; 12'd225: toneL = 32'd588; 
                12'd226: toneL = 32'd588; 12'd227: toneL = 32'd588; 
                12'd228: toneL = 32'd588; 12'd229: toneL = 32'd588; 
                12'd230: toneL = 32'd588; 12'd231: toneL = 32'd588; 
                12'd232: toneL = 32'd588; 12'd233: toneL = 32'd588; 
                12'd234: toneL = 32'd588; 12'd235: toneL = 32'd588; 
                12'd236: toneL = 32'd588; 12'd237: toneL = 32'd588; 
                12'd238: toneL = 32'd588; 12'd239: toneL = 32'd588; 
                12'd240: toneL = 32'd588; 12'd241: toneL = 32'd588; 
                12'd242: toneL = 32'd588; 12'd243: toneL = 32'd588; 
                12'd244: toneL = 32'd588; 12'd245: toneL = 32'd588; 
                12'd246: toneL = 32'd588; 12'd247: toneL = 32'd588; 
                12'd248: toneL = 32'd588; 12'd249: toneL = 32'd588; 
                12'd250: toneL = 32'd588; 12'd251: toneL = 32'd588; 
                12'd252: toneL = 32'd588; 12'd253: toneL = 32'd588; 
                12'd254: toneL = 32'd588; 12'd255: toneL = 32'd588;
                12'd256: toneL = 32'd588; 12'd257: toneL = 32'd588; 
                12'd258: toneL = 32'd588; 12'd259: toneL = 32'd588; 
                12'd260: toneL = 32'd588; 12'd261: toneL = 32'd588;
                12'd262: toneL = 32'd660; 12'd263: toneL = 32'd660;
                12'd264: toneL = 32'd524; 12'd265: toneL = 32'd524; 
                12'd266: toneL = 32'd524; 12'd267: toneL = 32'd524; 
                12'd268: toneL = 32'd524; 12'd269: toneL = 32'd524; 
                12'd270: toneL = 32'd524; 12'd271: toneL = 32'd524; 
                12'd272: toneL = 32'd524; 12'd273: toneL = 32'd524; 
                12'd274: toneL = 32'd524; 12'd275: toneL = 32'd524; 
                12'd276: toneL = 32'd524; 12'd277: toneL = 32'd524;
                12'd278: toneL = 32'd554; 12'd279: toneL = 32'd554;
                12'd280: toneL = 32'd588; 12'd281: toneL = 32'd588; 
                12'd282: toneL = 32'd588; 12'd283: toneL = 32'd588; 
                12'd284: toneL = 32'd588; 12'd285: toneL = 32'd588; 
                12'd286: toneL = 32'd588; 12'd287: toneL = 32'd588;
                12'd288: toneL = 32'd588; 12'd289: toneL = 32'd588; 
                12'd290: toneL = 32'd588; 12'd291: toneL = 32'd588; 
                12'd292: toneL = 32'd588; 12'd293: toneL = 32'd588;
                12'd294: toneL = 32'd660; 12'd295: toneL = 32'd660;
                12'd296: toneL = 32'd524; 12'd297: toneL = 32'd524; 
                12'd298: toneL = 32'd524; 12'd299: toneL = 32'd524; 
                12'd300: toneL = 32'd524; 12'd301: toneL = 32'd524; 
                12'd302: toneL = 32'd524; 12'd303: toneL = 32'd524; 
                12'd304: toneL = 32'd524; 12'd305: toneL = 32'd524; 
                12'd306: toneL = 32'd524; 12'd307: toneL = 32'd524; 
                12'd308: toneL = 32'd524; 12'd309: toneL = 32'd524; 
                12'd310: toneL = 32'd440; 12'd311: toneL = 32'd440;
                12'd312: toneL = 32'd392; 12'd313: toneL = 32'd392; 
                12'd314: toneL = 32'd392; 12'd315: toneL = 32'd392; 
                12'd316: toneL = 32'd392; 12'd317: toneL = 32'd392; 
                12'd318: toneL = 32'd392; 12'd319: toneL = 32'd392; 
                12'd320: toneL = 32'd392; 12'd321: toneL = 32'd392; 
                12'd322: toneL = 32'd392; 12'd323: toneL = 32'd392; 
                12'd324: toneL = 32'd392; 12'd325: toneL = 32'd392; 
                12'd326: toneL = 32'd392; 12'd327: toneL = 32'd392; 
                12'd328: toneL = 32'd330; 12'd329: toneL = 32'd330; 
                12'd330: toneL = 32'd330; 12'd331: toneL = 32'd330; 
                12'd332: toneL = 32'd330; 12'd333: toneL = 32'd330; 
                12'd334: toneL = 32'd330; 12'd335: toneL = 32'd330; 
                12'd336: toneL = 32'd330; 12'd337: toneL = 32'd330; 
                12'd338: toneL = 32'd330; 12'd339: toneL = 32'd330;
                12'd340: toneL = 32'd392; 12'd341: toneL = 32'd392; 
                12'd342: toneL = 32'd392; 12'd343: toneL = 32'd392; 
                12'd344: toneL = 32'd524; 12'd345: toneL = 32'd524; 
                12'd346: toneL = 32'd524; 12'd347: toneL = 32'd524; 
                12'd348: toneL = 32'd494; 12'd349: toneL = 32'd494; 
                12'd350: toneL = 32'd494; 12'd351: toneL = 32'd494; 
                12'd352: toneL = 32'd588; 12'd353: toneL = 32'd588; 
                12'd354: toneL = 32'd588; 12'd355: toneL = 32'd588; 
                12'd356: toneL = 32'd588; 12'd357: toneL = 32'd588; 
                12'd358: toneL = 32'd660; 12'd359: toneL = 32'd660;
                12'd360: toneL = 32'd524; 12'd361: toneL = 32'd524; 
                12'd362: toneL = 32'd524; 12'd363: toneL = 32'd524; 
                12'd364: toneL = 32'd524; 12'd365: toneL = 32'd524; 
                12'd366: toneL = 32'd524; 12'd367: toneL = 32'd524; 
                12'd368: toneL = 32'd524; 12'd369: toneL = 32'd524; 
                12'd370: toneL = 32'd524; 12'd371: toneL = 32'd524; 
                12'd372: toneL = 32'd524; 12'd373: toneL = 32'd524; 
                12'd374: toneL = 32'd554; 12'd375: toneL = 32'd554;
                12'd376: toneL = 32'd588; 12'd377: toneL = 32'd588; 
                12'd378: toneL = 32'd588; 12'd379: toneL = 32'd588; 
                12'd380: toneL = 32'd588; 12'd381: toneL = 32'd588; 
                12'd382: toneL = 32'd588; 12'd383: toneL = 32'd588; 
                12'd384: toneL = 32'd588; 12'd385: toneL = 32'd588; 
                12'd386: toneL = 32'd588; 12'd387: toneL = 32'd588; 
                12'd388: toneL = 32'd588; 12'd389: toneL = 32'd588; 
                12'd390: toneL = 32'd660; 12'd391: toneL = 32'd660;
                12'd392: toneL = 32'd524; 12'd393: toneL = 32'd524; 
                12'd394: toneL = 32'd524; 12'd395: toneL = 32'd524; 
                12'd396: toneL = 32'd524; 12'd397: toneL = 32'd524; 
                12'd398: toneL = 32'd524; 12'd399: toneL = 32'd524; 
                12'd400: toneL = 32'd524; 12'd401: toneL = 32'd524; 
                12'd402: toneL = 32'd524; 12'd403: toneL = 32'd524; 
                12'd404: toneL = 32'd524; 12'd405: toneL = 32'd524; 
                12'd406: toneL = 32'd440; 12'd407: toneL = 32'd440;
                12'd408: toneL = 32'd392; 12'd409: toneL = 32'd392; 
                12'd410: toneL = 32'd392; 12'd411: toneL = 32'd392; 
                12'd412: toneL = 32'd392; 12'd413: toneL = 32'd392; 
                12'd414: toneL = 32'd392; 12'd415: toneL = 32'd392; 
                12'd416: toneL = 32'd392; 12'd417: toneL = 32'd392; 
                12'd418: toneL = 32'd392; 12'd419: toneL = 32'd392; 
                12'd420: toneL = 32'd392; 12'd421: toneL = 32'd392; 
                12'd422: toneL = 32'd415; 12'd423: toneL = 32'd415;
                12'd424: toneL = 32'd440; 12'd425: toneL = 32'd440; 
                12'd426: toneL = 32'd440; 12'd427: toneL = 32'd440; 
                12'd428: toneL = 32'd440; 12'd429: toneL = 32'd440; 
                12'd430: toneL = 32'd440; 12'd431: toneL = 32'd440; 
                12'd432: toneL = 32'd440; 12'd433: toneL = 32'd440; 
                12'd434: toneL = 32'd440; 12'd435: toneL = 32'd440; 
                12'd436: toneL = 32'd466; 12'd437: toneL = 32'd466; 
                12'd438: toneL = 32'd466; 12'd439: toneL = 32'd466; 
                12'd440: toneL = 32'd494; 12'd441: toneL = 32'd494; 
                12'd442: toneL = 32'd494; 12'd443: toneL = 32'd494; 
                12'd444: toneL = 32'd494; 12'd445: toneL = 32'd494; 
                12'd446: toneL = 32'd494; 12'd447: toneL = 32'd494; 
                12'd448: toneL = 32'd494; 12'd449: toneL = 32'd494; 
                12'd450: toneL = 32'd494; 12'd451: toneL = 32'd494; 
                12'd452: toneL = 32'd392; 12'd453: toneL = 32'd392; 
                12'd454: toneL = 32'd392; 12'd455: toneL = 32'd392; 
                12'd456: toneL = 32'd524; 12'd457: toneL = 32'd524; 
                12'd458: toneL = 32'd524; 12'd459: toneL = 32'd524; 
                12'd460: toneL = 32'd524; 12'd461: toneL = 32'd524; 
                12'd462: toneL = 32'd524; 12'd463: toneL = 32'd524; 
                12'd464: toneL = 32'd494; 12'd465: toneL = 32'd494; 
                12'd466: toneL = 32'd494; 12'd467: toneL = 32'd494; 
                12'd468: toneL = 32'd494; 12'd469: toneL = 32'd494; 
                12'd470: toneL = 32'd524; 12'd471: toneL = 32'd524;
                12'd472: toneL = `sil; 12'd473: toneL = `sil; 
                12'd474: toneL = `sil; 12'd475: toneL = `sil; 
                12'd476: toneL = `sil; 12'd477: toneL = `sil; 
                12'd478: toneL = `sil; 12'd479: toneL = `sil; 
                12'd480: toneL = `sil; 12'd481: toneL = `sil; 
                12'd482: toneL = `sil; 12'd483: toneL = `sil; 
                12'd484: toneL = `sil; 12'd485: toneL = `sil; 
                12'd486: toneL = `sil; 12'd487: toneL = `sil; 
                12'd488: toneL = `sil; 12'd489: toneL = `sil; 
                12'd490: toneL = `sil; 12'd491: toneL = `sil; 
                12'd492: toneL = `sil; 12'd493: toneL = `sil; 
                12'd494: toneL = `sil; 12'd495: toneL = `sil; 
                12'd496: toneL = `sil; 12'd497: toneL = `sil; 
                12'd498: toneL = `sil; 12'd499: toneL = `sil; 
                12'd500: toneL = `sil; 12'd501: toneL = `sil; 
                12'd502: toneL = `sil; 12'd503: toneL = `sil; 
                12'd504: toneL = `sil; 12'd505: toneL = `sil; 
                12'd506: toneL = `sil; 12'd507: toneL = `sil; 
                12'd508: toneL = `sil; 12'd509: toneL = `sil; 
                12'd510: toneL = `sil; 12'd511: toneL = `sil; 
                12'd512: toneL = 32'd392; 12'd513: toneL = 32'd392; 
                12'd514: toneL = 32'd392; 12'd515: toneL = 32'd392; 
                12'd516: toneL = 32'd392; 12'd517: toneL = 32'd392; 
                12'd518: toneL = 32'd415; 12'd519: toneL = 32'd415;
                12'd520: toneL = 32'd440; 12'd521: toneL = 32'd440; 
                12'd522: toneL = 32'd440; 12'd523: toneL = 32'd440; 
                12'd524: toneL = 32'd440; 12'd525: toneL = 32'd440; 
                12'd526: toneL = 32'd440; 12'd527: toneL = 32'd440; 
                12'd528: toneL = 32'd440; 12'd529: toneL = 32'd440; 
                12'd530: toneL = 32'd440; 12'd531: toneL = 32'd440; 
                12'd532: toneL = 32'd440; 12'd533: toneL = 32'd440; 
                12'd534: toneL = 32'd440; 12'd535: toneL = 32'd440; 
                12'd536: toneL = 32'd440; 12'd537: toneL = 32'd440; 
                12'd538: toneL = 32'd440; 12'd539: toneL = 32'd440; 
                12'd540: toneL = 32'd440; 12'd541: toneL = 32'd440; 
                12'd542: toneL = 32'd440; 12'd543: toneL = 32'd440; 
                12'd544: toneL = 32'd440; 12'd545: toneL = 32'd440; 
                12'd546: toneL = 32'd440; 12'd547: toneL = 32'd440; 
                12'd548: toneL = 32'd440; 12'd549: toneL = 32'd440; 
                12'd550: toneL = 32'd440; 12'd551: toneL = 32'd440; 
                12'd552: toneL = 32'd440; 12'd553: toneL = 32'd440; 
                12'd554: toneL = 32'd440; 12'd555: toneL = 32'd440; 
                12'd556: toneL = 32'd440; 12'd557: toneL = 32'd440; 
                12'd558: toneL = 32'd392; 12'd559: toneL = 32'd392;
                12'd560: toneL = 32'd440; 12'd561: toneL = 32'd440; 
                12'd562: toneL = 32'd440; 12'd563: toneL = 32'd440; 
                12'd564: toneL = 32'd440; 12'd565: toneL = 32'd440; 
                12'd566: toneL = 32'd392; 12'd567: toneL = 32'd392;
                12'd568: toneL = 32'd440; 12'd569: toneL = 32'd440; 
                12'd570: toneL = 32'd440; 12'd571: toneL = 32'd440; 
                12'd572: toneL = 32'd440; 12'd573: toneL = 32'd440;
                12'd574: toneL = 32'd392; 12'd575: toneL = 32'd392;
                12'd576: toneL = 32'd330; 12'd577: toneL = 32'd330; 
                12'd578: toneL = 32'd330; 12'd579: toneL = 32'd330; 
                12'd580: toneL = 32'd330; 12'd581: toneL = 32'd330; 
                12'd582: toneL = 32'd262; 12'd583: toneL = 32'd262;
                12'd584: toneL = 32'd440; 12'd585: toneL = 32'd440; 
                12'd586: toneL = 32'd440; 12'd587: toneL = 32'd440; 
                12'd588: toneL = 32'd440; 12'd589: toneL = 32'd440; 
                12'd590: toneL = 32'd440; 12'd591: toneL = 32'd440; 
                12'd592: toneL = 32'd440; 12'd593: toneL = 32'd440; 
                12'd594: toneL = 32'd440; 12'd595: toneL = 32'd440; 
                12'd596: toneL = 32'd440; 12'd597: toneL = 32'd440; 
                12'd598: toneL = 32'd440; 12'd599: toneL = 32'd440; 
                12'd600: toneL = 32'd440; 12'd601: toneL = 32'd440; 
                12'd602: toneL = 32'd440; 12'd603: toneL = 32'd440; 
                12'd604: toneL = 32'd440; 12'd605: toneL = 32'd440; 
                12'd606: toneL = 32'd440; 12'd607: toneL = 32'd440; 
                12'd608: toneL = 32'd440; 12'd609: toneL = 32'd440; 
                12'd610: toneL = 32'd440; 12'd611: toneL = 32'd440; 
                12'd612: toneL = 32'd440; 12'd613: toneL = 32'd440; 
                12'd614: toneL = 32'd440; 12'd615: toneL = 32'd440; 
                12'd616: toneL = 32'd440; 12'd617: toneL = 32'd440; 
                12'd618: toneL = 32'd440; 12'd619: toneL = 32'd440; 
                12'd620: toneL = 32'd440; 12'd621: toneL = 32'd440; 
                12'd622: toneL = 32'd440; 12'd623: toneL = 32'd440; 
                12'd624: toneL = 32'd440; 12'd625: toneL = 32'd440; 
                12'd626: toneL = 32'd440; 12'd627: toneL = 32'd440; 
                12'd628: toneL = 32'd440; 12'd629: toneL = 32'd440; 
                12'd630: toneL = 32'd440; 12'd631: toneL = 32'd440; 
                12'd632: toneL = 32'd440; 12'd633: toneL = 32'd440; 
                12'd634: toneL = 32'd440; 12'd635: toneL = 32'd440; 
                12'd636: toneL = 32'd440; 12'd637: toneL = 32'd440; 
                12'd638: toneL = 32'd440; 12'd639: toneL = 32'd440; 
                12'd640: toneL = 32'd524; 12'd641: toneL = 32'd524; 
                12'd642: toneL = 32'd524; 12'd643: toneL = 32'd524; 
                12'd644: toneL = 32'd524; 12'd645: toneL = 32'd524; 
                12'd646: toneL = 32'd554; 12'd647: toneL = 32'd554;
                12'd648: toneL = 32'd588; 12'd649: toneL = 32'd588; 
                12'd650: toneL = 32'd588; 12'd651: toneL = 32'd588; 
                12'd652: toneL = 32'd588; 12'd653: toneL = 32'd588; 
                12'd654: toneL = 32'd588; 12'd655: toneL = 32'd588; 
                12'd656: toneL = 32'd588; 12'd657: toneL = 32'd588; 
                12'd658: toneL = 32'd588; 12'd659: toneL = 32'd588; 
                12'd660: toneL = 32'd588; 12'd661: toneL = 32'd588; 
                12'd662: toneL = 32'd588; 12'd663: toneL = 32'd588; 
                12'd664: toneL = 32'd588; 12'd665: toneL = 32'd588; 
                12'd666: toneL = 32'd588; 12'd667: toneL = 32'd588; 
                12'd668: toneL = 32'd588; 12'd669: toneL = 32'd588; 
                12'd670: toneL = 32'd588; 12'd671: toneL = 32'd588; 
                12'd672: toneL = 32'd588; 12'd673: toneL = 32'd588; 
                12'd674: toneL = 32'd588; 12'd675: toneL = 32'd588; 
                12'd676: toneL = 32'd588; 12'd677: toneL = 32'd588; 
                12'd678: toneL = 32'd588; 12'd679: toneL = 32'd588; 
                12'd680: toneL = 32'd588; 12'd681: toneL = 32'd588; 
                12'd682: toneL = 32'd588; 12'd683: toneL = 32'd588; 
                12'd684: toneL = 32'd588; 12'd685: toneL = 32'd588; 
                12'd686: toneL = 32'd660; 12'd687: toneL = 32'd660;
                12'd688: toneL = 32'd588; 12'd689: toneL = 32'd588; 
                12'd690: toneL = 32'd588; 12'd691: toneL = 32'd588; 
                12'd692: toneL = 32'd588; 12'd693: toneL = 32'd588; 
                12'd694: toneL = 32'd660; 12'd695: toneL = 32'd660;
                12'd696: toneL = 32'd588; 12'd697: toneL = 32'd588; 
                12'd698: toneL = 32'd588; 12'd699: toneL = 32'd588; 
                12'd700: toneL = 32'd588; 12'd701: toneL = 32'd588; 
                12'd702: toneL = 32'd524; 12'd703: toneL = 32'd524; 
                12'd704: toneL = 32'd524; 12'd705: toneL = 32'd524; 
                12'd706: toneL = 32'd415; 12'd707: toneL = 32'd415;
                12'd708: toneL = 32'd349; 12'd709: toneL = 32'd349;
                12'd710: toneL = 32'd588; 12'd711: toneL = 32'd588; 
                12'd712: toneL = 32'd588; 12'd713: toneL = 32'd588; 
                12'd714: toneL = 32'd588; 12'd715: toneL = 32'd588; 
                12'd716: toneL = 32'd588; 12'd717: toneL = 32'd588; 
                12'd718: toneL = 32'd588; 12'd719: toneL = 32'd588; 
                12'd720: toneL = 32'd588; 12'd721: toneL = 32'd588; 
                12'd722: toneL = 32'd588; 12'd723: toneL = 32'd588; 
                12'd724: toneL = 32'd588; 12'd725: toneL = 32'd588; 
                12'd726: toneL = 32'd588; 12'd727: toneL = 32'd588; 
                12'd728: toneL = 32'd588; 12'd729: toneL = 32'd588; 
                12'd730: toneL = 32'd588; 12'd731: toneL = 32'd588; 
                12'd732: toneL = 32'd588; 12'd733: toneL = 32'd588; 
                12'd734: toneL = 32'd588; 12'd735: toneL = 32'd588; 
                12'd736: toneL = 32'd588; 12'd737: toneL = 32'd588; 
                12'd738: toneL = 32'd588; 12'd739: toneL = 32'd588; 
                12'd740: toneL = 32'd588; 12'd741: toneL = 32'd588; 
                12'd742: toneL = 32'd588; 12'd743: toneL = 32'd588; 
                12'd744: toneL = 32'd588; 12'd745: toneL = 32'd588; 
                12'd746: toneL = 32'd588; 12'd747: toneL = 32'd588; 
                12'd748: toneL = 32'd588; 12'd749: toneL = 32'd588; 
                12'd750: toneL = 32'd588; 12'd751: toneL = 32'd588; 
                12'd752: toneL = 32'd588; 12'd753: toneL = 32'd588; 
                12'd754: toneL = 32'd588; 12'd755: toneL = 32'd588; 
                12'd756: toneL = 32'd588; 12'd757: toneL = 32'd588; 
                12'd758: toneL = 32'd588; 12'd759: toneL = 32'd588; 
                12'd760: toneL = 32'd588; 12'd761: toneL = 32'd588; 
                12'd762: toneL = 32'd588; 12'd763: toneL = 32'd588; 
                12'd764: toneL = 32'd588; 12'd765: toneL = 32'd588; 
                12'd766: toneL = 32'd588; 12'd767: toneL = 32'd588; 
                12'd768: toneL = 32'd588; 12'd769: toneL = 32'd588; 
                12'd770: toneL = 32'd588; 12'd771: toneL = 32'd588; 
                12'd772: toneL = 32'd588; 12'd773: toneL = 32'd588; 
                12'd774: toneL = 32'd660; 12'd775: toneL = 32'd660;
                12'd776: toneL = 32'd524; 12'd777: toneL = 32'd524; 
                12'd778: toneL = 32'd524; 12'd779: toneL = 32'd524; 
                12'd780: toneL = 32'd524; 12'd781: toneL = 32'd524; 
                12'd782: toneL = 32'd524; 12'd783: toneL = 32'd524; 
                12'd784: toneL = 32'd524; 12'd785: toneL = 32'd524; 
                12'd786: toneL = 32'd524; 12'd787: toneL = 32'd524; 
                12'd788: toneL = 32'd524; 12'd789: toneL = 32'd524;
                12'd790: toneL = 32'd554; 12'd791: toneL = 32'd554;
                12'd792: toneL = 32'd588; 12'd793: toneL = 32'd588; 
                12'd794: toneL = 32'd588; 12'd795: toneL = 32'd588; 
                12'd796: toneL = 32'd588; 12'd797: toneL = 32'd588; 
                12'd798: toneL = 32'd588; 12'd799: toneL = 32'd588; 
                12'd800: toneL = 32'd588; 12'd801: toneL = 32'd588; 
                12'd802: toneL = 32'd588; 12'd803: toneL = 32'd588; 
                12'd804: toneL = 32'd588; 12'd805: toneL = 32'd588; 
                12'd806: toneL = 32'd660; 12'd807: toneL = 32'd660;
                12'd808: toneL = 32'd524; 12'd809: toneL = 32'd524; 
                12'd810: toneL = 32'd524; 12'd811: toneL = 32'd524; 
                12'd812: toneL = 32'd524; 12'd813: toneL = 32'd524; 
                12'd814: toneL = 32'd524; 12'd815: toneL = 32'd524; 
                12'd816: toneL = 32'd524; 12'd817: toneL = 32'd524; 
                12'd818: toneL = 32'd524; 12'd819: toneL = 32'd524; 
                12'd820: toneL = 32'd524; 12'd821: toneL = 32'd524; 
                12'd822: toneL = 32'd440; 12'd823: toneL = 32'd440;
                12'd824: toneL = 32'd392; 12'd825: toneL = 32'd392; 
                12'd826: toneL = 32'd392; 12'd827: toneL = 32'd392; 
                12'd828: toneL = 32'd392; 12'd829: toneL = 32'd392; 
                12'd830: toneL = 32'd392; 12'd831: toneL = 32'd392; 
                12'd832: toneL = 32'd392; 12'd833: toneL = 32'd392; 
                12'd834: toneL = 32'd392; 12'd835: toneL = 32'd392; 
                12'd836: toneL = 32'd392; 12'd837: toneL = 32'd392; 
                12'd838: toneL = 32'd392; 12'd839: toneL = 32'd392; 
                12'd840: toneL = 32'd330; 12'd841: toneL = 32'd330; 
                12'd842: toneL = 32'd330; 12'd843: toneL = 32'd330; 
                12'd844: toneL = 32'd330; 12'd845: toneL = 32'd330; 
                12'd846: toneL = 32'd330; 12'd847: toneL = 32'd330; 
                12'd848: toneL = 32'd330; 12'd849: toneL = 32'd330; 
                12'd850: toneL = 32'd330; 12'd851: toneL = 32'd330; 
                12'd852: toneL = 32'd392; 12'd853: toneL = 32'd392; 
                12'd854: toneL = 32'd392; 12'd855: toneL = 32'd392; 
                12'd856: toneL = 32'd524; 12'd857: toneL = 32'd524; 
                12'd858: toneL = 32'd524; 12'd859: toneL = 32'd524; 
                12'd860: toneL = 32'd494; 12'd861: toneL = 32'd494; 
                12'd862: toneL = 32'd494; 12'd863: toneL = 32'd494; 
                12'd864: toneL = 32'd588; 12'd865: toneL = 32'd588; 
                12'd866: toneL = 32'd588; 12'd867: toneL = 32'd588; 
                12'd868: toneL = 32'd588; 12'd869: toneL = 32'd588; 
                12'd870: toneL = 32'd660; 12'd871: toneL = 32'd660;
                12'd872: toneL = 32'd524; 12'd873: toneL = 32'd524; 
                12'd874: toneL = 32'd524; 12'd875: toneL = 32'd524; 
                12'd876: toneL = 32'd524; 12'd877: toneL = 32'd524; 
                12'd878: toneL = 32'd524; 12'd879: toneL = 32'd524; 
                12'd880: toneL = 32'd524; 12'd881: toneL = 32'd524; 
                12'd882: toneL = 32'd524; 12'd883: toneL = 32'd524; 
                12'd884: toneL = 32'd524; 12'd885: toneL = 32'd524; 
                12'd886: toneL = 32'd554; 12'd887: toneL = 32'd554;
                12'd888: toneL = 32'd588; 12'd889: toneL = 32'd588; 
                12'd890: toneL = 32'd588; 12'd891: toneL = 32'd588; 
                12'd892: toneL = 32'd588; 12'd893: toneL = 32'd588; 
                12'd894: toneL = 32'd588; 12'd895: toneL = 32'd588; 
                12'd896: toneL = 32'd588; 12'd897: toneL = 32'd588; 
                12'd898: toneL = 32'd588; 12'd899: toneL = 32'd588; 
                12'd900: toneL = 32'd588; 12'd901: toneL = 32'd588; 
                12'd902: toneL = 32'd660; 12'd903: toneL = 32'd660;
                12'd904: toneL = 32'd524; 12'd905: toneL = 32'd524; 
                12'd906: toneL = 32'd524; 12'd907: toneL = 32'd524; 
                12'd908: toneL = 32'd524; 12'd909: toneL = 32'd524; 
                12'd910: toneL = 32'd524; 12'd911: toneL = 32'd524; 
                12'd912: toneL = 32'd524; 12'd913: toneL = 32'd524; 
                12'd914: toneL = 32'd524; 12'd915: toneL = 32'd524; 
                12'd916: toneL = 32'd524; 12'd917: toneL = `sil; 
                12'd918: toneL = 32'd440; 12'd919: toneL = 32'd440;
                12'd920: toneL = 32'd392; 12'd921: toneL = 32'd392; 
                12'd922: toneL = 32'd392; 12'd923: toneL = 32'd392; 
                12'd924: toneL = 32'd392; 12'd925: toneL = 32'd392; 
                12'd926: toneL = 32'd392; 12'd927: toneL = 32'd392; 
                12'd928: toneL = 32'd392; 12'd929: toneL = 32'd392; 
                12'd930: toneL = 32'd392; 12'd931: toneL = 32'd392; 
                12'd932: toneL = 32'd392; 12'd933: toneL = 32'd392;
                12'd934: toneL = 32'd415; 12'd935: toneL = 32'd415;
                12'd936: toneL = 32'd440; 12'd937: toneL = 32'd440; 
                12'd938: toneL = 32'd440; 12'd939: toneL = 32'd440; 
                12'd940: toneL = 32'd440; 12'd941: toneL = 32'd440; 
                12'd942: toneL = 32'd440; 12'd943: toneL = 32'd440; 
                12'd944: toneL = 32'd440; 12'd945: toneL = 32'd440; 
                12'd946: toneL = 32'd440; 12'd947: toneL = 32'd440; 
                12'd948: toneL = 32'd466; 12'd949: toneL = 32'd466; 
                12'd950: toneL = 32'd466; 12'd951: toneL = 32'd466; 
                12'd952: toneL = 32'd494; 12'd953: toneL = 32'd494; 
                12'd954: toneL = 32'd494; 12'd955: toneL = 32'd494; 
                12'd956: toneL = 32'd494; 12'd957: toneL = 32'd494; 
                12'd958: toneL = 32'd494; 12'd959: toneL = 32'd494; 
                12'd960: toneL = 32'd494; 12'd961: toneL = 32'd494; 
                12'd962: toneL = 32'd494; 12'd963: toneL = 32'd494; 
                12'd964: toneL = 32'd392; 12'd965: toneL = 32'd392; 
                12'd966: toneL = 32'd392; 12'd967: toneL = 32'd392; 
                12'd968: toneL = 32'd524; 12'd969: toneL = 32'd524; 
                12'd970: toneL = 32'd524; 12'd971: toneL = 32'd524; 
                12'd972: toneL = 32'd524; 12'd973: toneL = 32'd524; 
                12'd974: toneL = 32'd524; 12'd975: toneL = 32'd524; 
                12'd976: toneL = 32'd494; 12'd977: toneL = 32'd494; 
                12'd978: toneL = 32'd494; 12'd979: toneL = 32'd494; 
                12'd980: toneL = 32'd494; 12'd981: toneL = 32'd494; 
                12'd982: toneL = 32'd524; 12'd983: toneL = 32'd524;
                12'd984: toneL = `sil; 12'd985: toneL = `sil; 
                12'd986: toneL = `sil; 12'd987: toneL = `sil; 
                12'd988: toneL = `sil; 12'd989: toneL = `sil; 
                12'd990: toneL = `sil; 12'd991: toneL = `sil; 
                12'd992: toneL = `sil; 12'd993: toneL = `sil; 
                12'd994: toneL = `sil; 12'd995: toneL = `sil; 
                12'd996: toneL = `sil; 12'd997: toneL = `sil; 
                12'd998: toneL = `sil; 12'd999: toneL = `sil; 
                12'd1000: toneL = `sil; 12'd1001: toneL = `sil; 
                12'd1002: toneL = `sil; 12'd1003: toneL = `sil; 
                12'd1004: toneL = `sil; 12'd1005: toneL = `sil; 
                12'd1006: toneL = `sil; 12'd1007: toneL = `sil; 
                12'd1008: toneL = `sil; 12'd1009: toneL = `sil; 
                12'd1010: toneL = `sil; 12'd1011: toneL = `sil; 
                12'd1012: toneL = `sil; 12'd1013: toneL = `sil; 
                12'd1014: toneL = `sil; 12'd1015: toneL = `sil; 
                12'd1016: toneL = `sil; 12'd1017: toneL = `sil; 
                12'd1018: toneL = `sil; 12'd1019: toneL = `sil; 
                12'd1020: toneL = `sil; 12'd1021: toneL = `sil; 
                12'd1022: toneL = `sil; 12'd1023: toneL = `sil; 



                default : toneL = `sil;
            endcase
        end
    end
endmodule